/* AUTHOR
* David Little
*/

`ifndef CHRONO_H_
`define CHRONO_H_

`include "globals.vh"



parameter   ROUND_DELAY = SECOND,
            SUCCESS_DELAY = MILLI_SECOND * 450,
            FAILURE_DELAY = SECOND,
            RECITE_MOVES_DELAY = SECOND,
            GAME_MOVE_LIGHT_DELAY = MILLI_SECOND * 202,
            GAME_MOVE_DARK_DELAY = MILLI_SECOND * 650,
            PLAYER_DO_MOVES_DELAY = MILLI_SECOND * 250;
    


`endif